//: version "2.1"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "lab5a.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg w3;    //: /sn:0 {0}(768,355)(768,465)(462,465){1}
//: {2}(460,463)(460,357){3}
//: {4}(460,467)(460,486){5}
reg w10;    //: /sn:0 {0}(230,216)(274,216){1}
//: {2}(278,216)(357,216){3}
//: {4}(361,216)(582,216){5}
//: {6}(586,216)(620,216){7}
//: {8}(624,216)(881,216)(881,162){9}
//: {10}(622,218)(622,264)(644,264){11}
//: {12}(584,218)(584,325)(698,325){13}
//: {14}(359,218)(359,264)(390,264){15}
//: {16}(276,218)(276,332)(311,332){17}
reg w11;    //: /sn:0 {0}(698,293)(631,293)(631,405)(344,405){1}
//: {2}(342,403)(342,295)(390,295){3}
//: {4}(340,405)(232,405){5}
wire w16;    //: /sn:0 {0}(552,325)(531,325){1}
wire w4;    //: /sn:0 {0}(390,332)(327,332){1}
wire w1;    //: /sn:0 {0}(884,141)(884,122){1}
wire w8;    //: /sn:0 {0}(839,323)(854,323){1}
wire w15;    //: /sn:0 {0}(531,269)(644,269){1}
wire w5;    //: /sn:0 {0}(665,267)(698,267){1}
wire w9;    //: /sn:0 {0}(839,267)(886,267)(886,162){1}
//: enddecls

  //: comment g4 @(266,383) /sn:0
  //: /line:"CLK"
  //: /end
  //: joint g8 (w3) @(460, 465) /w:[ 1 2 -1 4 ]
  //: SWITCH X (w10) @(213,216) /w:[ 0 ] /st:1 /dn:0
  _GGAND2 #(6) g16 (.I0(!w10), .I1(w9), .Z(w1));   //: @(884,151) /sn:0 /R:1 /w:[ 9 1 0 ]
  //: joint g18 (w10) @(584, 216) /w:[ 6 -1 5 12 ]
  //: LED Z (w1) @(884,115) /w:[ 1 ] /type:0
  //: SWITCH RESET (w3) @(460,500) /sn:0 /R:1 /w:[ 5 ] /st:1 /dn:0
  JKFlipFlop JK1 (.CLK(w11), .K(w4), .J(w10), .Reset(w3), .Qinv(w16), .Q(w15));   //: @(391, 241) /sz:(139, 115) /p:[ Li0>3 Li1>0 Li2>15 Bi0>3 Ro0<1 Ro1<0 ]
  //: joint g12 (w10) @(276, 216) /w:[ 2 -1 1 16 ]
  _GGAND2 #(6) g14 (.I0(!w10), .I1(w15), .Z(w5));   //: @(655,267) /sn:0 /w:[ 11 1 0 ]
  //: joint g11 (w10) @(359, 216) /w:[ 4 -1 3 14 ]
  //: joint g5 (w11) @(342, 405) /w:[ 1 2 4 -1 ]
  JKFlipFlop JK0 (.J(w5), .K(w10), .CLK(w11), .Reset(w3), .Q(w9), .Qinv(w8));   //: @(699, 239) /sz:(139, 115) /sn:0 /p:[ Li0>1 Li1>13 Li2>0 Bi0>0 Ro0<0 Ro1<0 ]
  //: SWITCH CLK (w11) @(215,405) /w:[ 5 ] /st:1 /dn:1
  //: joint g15 (w10) @(622, 216) /w:[ 8 -1 7 10 ]
  _GGNBUF #(2) g13 (.I(w10), .Z(w4));   //: @(317,332) /sn:0 /w:[ 17 1 ]

endmodule
//: /netlistEnd

//: /netlistBegin JKFlipFlop
module JKFlipFlop(K, J, Reset, CLK, Qinv, Q);
//: interface  /sz:(139, 115) /bd:[ Li0>J(23/115) Li1>K(86/115) Li2>CLK(54/115) Bi0>Reset(69/139) Ro0<Q(28/115) Ro1<Qinv(84/115) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
output Q;    //: /sn:0 {0}(299,274)(284,274)(284,315)(682,315)(682,220){1}
//: {2}(684,218)(696,218)(696,217)(706,217){3}
//: {4}(680,218)(652,218){5}
//: {6}(648,218)(629,218){7}
//: {8}(650,220)(650,257)(592,257)(592,265)(608,265){9}
input K;    //: /sn:0 {0}(180,279)(299,279){1}
input J;    //: /sn:0 {0}(185,205)(301,205){1}
output Qinv;    //: /sn:0 {0}(710,270)(672,270){1}
//: {2}(670,268)(670,178)(281,178)(281,210)(301,210){3}
//: {4}(668,270)(661,270){5}
//: {6}(659,268)(659,236)(594,236)(594,220)(608,220){7}
//: {8}(657,270)(629,270){9}
input Reset;    //: /sn:0 {0}(589,311)(589,310){1}
//: {2}(589,306)(589,275)(608,275){3}
//: {4}(587,308)(469,308){5}
//: {6}(465,308)(387,308)(387,284)(398,284){7}
//: {8}(467,310)(467,358){9}
input CLK;    //: /sn:0 {0}(197,335)(291,335){1}
//: {2}(295,335)(305,335){3}
//: {4}(293,333)(293,330)(305,330){5}
//: {6}(293,337)(293,347)(278,347)(278,269)(290,269){7}
//: {8}(294,269)(299,269){9}
//: {10}(292,267)(292,215)(301,215){11}
wire w13;    //: /sn:0 {0}(534,270)(608,270){1}
wire w7;    //: /sn:0 {0}(419,279)(448,279){1}
//: {2}(452,279)(498,279)(498,272)(513,272){3}
//: {4}(450,277)(450,236)(381,236)(381,214)(391,214){5}
wire w8;    //: /sn:0 {0}(398,279)(383,279)(383,249)(434,249)(434,214){1}
//: {2}(436,212)(511,212){3}
//: {4}(432,212)(412,212){5}
wire w14;    //: /sn:0 {0}(532,215)(608,215){1}
wire w2;    //: /sn:0 {0}(322,210)(376,210)(376,209)(391,209){1}
wire w5;    //: /sn:0 {0}(320,274)(398,274){1}
wire w26;    //: /sn:0 {0}(511,217)(488,217)(488,265){1}
//: {2}(490,267)(513,267){3}
//: {4}(488,269)(488,333)(326,333){5}
//: enddecls

  _GGNAND2 #(4) g8 (.I0(CLK), .I1(CLK), .Z(w26));   //: @(316,333) /sn:0 /w:[ 5 3 5 ]
  _GGNAND2 #(4) g4 (.I0(w8), .I1(w26), .Z(w14));   //: @(522,215) /sn:0 /w:[ 3 0 0 ]
  _GGNAND3 #(6) g3 (.I0(w5), .I1(w8), .I2(Reset), .Z(w7));   //: @(409,279) /sn:0 /w:[ 1 0 7 0 ]
  //: joint g16 (CLK) @(292, 269) /w:[ 8 10 7 -1 ]
  //: joint g17 (Reset) @(467, 308) /w:[ 5 -1 6 8 ]
  _GGNAND2 #(4) g2 (.I0(w2), .I1(w7), .Z(w8));   //: @(402,212) /sn:0 /w:[ 1 5 5 ]
  //: joint g23 (Q) @(650, 218) /w:[ 5 -1 6 8 ]
  _GGNAND3 #(6) g1 (.I0(CLK), .I1(Q), .I2(K), .Z(w5));   //: @(310,274) /sn:0 /w:[ 9 0 1 0 ]
  //: joint g24 (Qinv) @(670, 270) /w:[ 1 2 4 -1 ]
  //: joint g18 (Reset) @(589, 308) /w:[ -1 2 4 1 ]
  //: IN g10 (K) @(178,279) /sn:0 /w:[ 0 ]
  //: joint g25 (Q) @(682, 218) /w:[ 2 -1 4 1 ]
  _GGNAND2 #(4) g6 (.I0(w14), .I1(Qinv), .Z(Q));   //: @(619,218) /sn:0 /w:[ 1 7 7 ]
  //: IN g9 (J) @(183,205) /sn:0 /w:[ 0 ]
  _GGNAND3 #(6) g7 (.I0(Q), .I1(w13), .I2(Reset), .Z(Qinv));   //: @(619,270) /sn:0 /w:[ 9 1 3 9 ]
  //: joint g22 (Qinv) @(659, 270) /w:[ 5 6 8 -1 ]
  //: IN g12 (Reset) @(467,360) /sn:0 /R:1 /w:[ 9 ]
  //: IN g11 (CLK) @(195,335) /sn:0 /w:[ 0 ]
  //: OUT g14 (Qinv) @(707,270) /sn:0 /w:[ 0 ]
  _GGNAND2 #(4) g5 (.I0(w26), .I1(w7), .Z(w13));   //: @(524,270) /sn:0 /w:[ 3 3 0 ]
  //: joint g19 (w26) @(488, 267) /w:[ 2 1 -1 4 ]
  //: joint g21 (w8) @(434, 212) /w:[ 2 -1 4 1 ]
  //: joint g20 (w7) @(450, 279) /w:[ 2 4 1 -1 ]
  //: joint g15 (CLK) @(293, 335) /w:[ 2 4 1 6 ]
  _GGNAND3 #(6) g0 (.I0(J), .I1(Qinv), .I2(CLK), .Z(w2));   //: @(312,210) /sn:0 /w:[ 1 3 11 0 ]
  //: OUT g13 (Q) @(703,217) /sn:0 /w:[ 3 ]

endmodule
//: /netlistEnd

