//: version "2.1"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "lab5a.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg w0;    //: /sn:0 {0}(473,302)(371,302){1}
//: {2}(367,302)(216,302){3}
//: {4}(369,304)(369,316)(369,316)(369,326){5}
reg w17;    //: /sn:0 {0}(1040,398)(1040,570)(799,570){1}
//: {2}(797,568)(797,395){3}
//: {4}(795,570)(545,570){5}
//: {6}(543,568)(543,394){7}
//: {8}(543,572)(543,589){9}
reg w2;    //: /sn:0 {0}(970,336)(935,336)(935,535)(686,535){1}
//: {2}(684,533)(684,333)(727,333){3}
//: {4}(682,535)(460,535){5}
//: {6}(458,533)(458,332)(473,332){7}
//: {8}(456,535)(322,535){9}
wire w6;    //: /sn:0 {0}(1111,310)(1121,310)(1121,263)(907,263)(907,156){1}
wire w4;    //: /sn:0 {0}(614,362)(727,362){1}
wire [2:0] w3;    //: /sn:0 {0}(#:897,150)(897,96){1}
wire w10;    //: /sn:0 {0}(868,363)(970,363){1}
wire w1;    //: /sn:0 {0}(369,342)(369,364)(473,364){1}
wire w11;    //: /sn:0 {0}(970,307)(899,307){1}
//: {2}(897,305)(897,156){3}
//: {4}(895,307)(868,307){5}
wire Q2;    //: /sn:0 {0}(614,305)(649,305){1}
//: {2}(653,305)(727,305){3}
//: {4}(651,303)(651,266)(887,266)(887,156){5}
wire w15;    //: /sn:0 {0}(1111,366)(1126,366){1}
//: enddecls

  JKFlipFlop A0 (.J(w0), .K(w1), .CLK(w2), .Reset(w17), .Q(Q2), .Qinv(w4));   //: @(474, 278) /sz:(139, 115) /p:[ Li0>0 Li1>1 Li2>7 Bi0>7 Ro0<0 Ro1<0 ]
  //: joint g8 (w17) @(797, 570) /w:[ 1 2 4 -1 ]
  //: joint g4 (w0) @(369, 302) /w:[ 1 -1 2 4 ]
  //: SWITCH X (w0) @(199,302) /w:[ 3 ] /st:0 /dn:0
  _GGNBUF #(2) g3 (.I(w0), .Z(w1));   //: @(369,332) /sn:0 /R:3 /w:[ 5 0 ]
  //: joint g10 (w2) @(684, 535) /w:[ 1 2 4 -1 ]
  JKFlipFlop A2 (.J(w11), .K(w10), .CLK(w2), .Reset(w17), .Q(w6), .Qinv(w15));   //: @(971, 282) /sz:(139, 115) /p:[ Li0>0 Li1>1 Li2>0 Bi0>0 Ro0<0 Ro1<0 ]
  //: SWITCH RESET (w17) @(543,603) /R:1 /w:[ 9 ] /st:0 /dn:0
  assign w3 = {w6, w11, Q2}; //: CONCAT g6  @(897,151) /sn:0 /R:1 /w:[ 0 1 3 5 ] /dr:1 /tp:0 /drp:1
  //: joint g9 (w2) @(458, 535) /w:[ 5 6 8 -1 ]
  //: joint g7 (w17) @(543, 570) /w:[ 5 6 -1 8 ]
  //: joint g12 (w11) @(897, 307) /w:[ 1 2 4 -1 ]
  //: joint g11 (Q2) @(651, 305) /w:[ 2 4 1 -1 ]
  //: LED g5 (w3) @(897,89) /sn:0 /w:[ 1 ] /type:3
  //: SWITCH CLK (w2) @(305,535) /w:[ 9 ] /st:0 /dn:0
  JKFlipFlop A1 (.J(Q2), .K(w4), .CLK(w2), .Reset(w17), .Q(w11), .Qinv(w10));   //: @(728, 279) /sz:(139, 115) /p:[ Li0>3 Li1>1 Li2>3 Bi0>3 Ro0<5 Ro1<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin JKFlipFlop
module JKFlipFlop(K, J, Reset, Qinv, CLK, Q);
//: interface  /sz:(139, 115) /bd:[ Li0>CLK(54/115) Li1>K(86/115) Li2>J(23/115) Bi0>Reset(69/139) Ro0<Qinv(84/115) Ro1<Q(28/115) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
output Q;    //: /sn:0 {0}(299,274)(284,274)(284,315)(682,315)(682,220){1}
//: {2}(684,218)(696,218)(696,217)(706,217){3}
//: {4}(680,218)(652,218){5}
//: {6}(648,218)(629,218){7}
//: {8}(650,220)(650,257)(592,257)(592,265)(608,265){9}
input K;    //: /sn:0 {0}(180,279)(299,279){1}
output Qinv;    //: /sn:0 {0}(710,270)(672,270){1}
//: {2}(670,268)(670,178)(281,178)(281,210)(301,210){3}
//: {4}(668,270)(661,270){5}
//: {6}(659,268)(659,236)(594,236)(594,220)(608,220){7}
//: {8}(657,270)(629,270){9}
input J;    //: /sn:0 {0}(185,205)(301,205){1}
input Reset;    //: /sn:0 {0}(589,311)(589,310){1}
//: {2}(589,306)(589,275)(608,275){3}
//: {4}(587,308)(469,308){5}
//: {6}(465,308)(387,308)(387,284)(398,284){7}
//: {8}(467,310)(467,358){9}
input CLK;    //: /sn:0 {0}(197,335)(291,335){1}
//: {2}(295,335)(305,335){3}
//: {4}(293,333)(293,330)(305,330){5}
//: {6}(293,337)(293,347)(278,347)(278,269)(290,269){7}
//: {8}(294,269)(299,269){9}
//: {10}(292,267)(292,215)(301,215){11}
wire w13;    //: /sn:0 {0}(534,270)(608,270){1}
wire w7;    //: /sn:0 {0}(419,279)(448,279){1}
//: {2}(452,279)(498,279)(498,272)(513,272){3}
//: {4}(450,277)(450,236)(381,236)(381,214)(391,214){5}
wire w8;    //: /sn:0 {0}(398,279)(383,279)(383,249)(434,249)(434,214){1}
//: {2}(436,212)(511,212){3}
//: {4}(432,212)(412,212){5}
wire w14;    //: /sn:0 {0}(532,215)(608,215){1}
wire w2;    //: /sn:0 {0}(322,210)(376,210)(376,209)(391,209){1}
wire w5;    //: /sn:0 {0}(320,274)(398,274){1}
wire w26;    //: /sn:0 {0}(511,217)(488,217)(488,265){1}
//: {2}(490,267)(513,267){3}
//: {4}(488,269)(488,333)(326,333){5}
//: enddecls

  _GGNAND2 #(4) g4 (.I0(w8), .I1(w26), .Z(w14));   //: @(522,215) /sn:0 /w:[ 3 0 0 ]
  _GGNAND2 #(4) g8 (.I0(CLK), .I1(CLK), .Z(w26));   //: @(316,333) /sn:0 /w:[ 5 3 5 ]
  //: joint g16 (CLK) @(292, 269) /w:[ 8 10 7 -1 ]
  _GGNAND3 #(6) g3 (.I0(w5), .I1(w8), .I2(Reset), .Z(w7));   //: @(409,279) /sn:0 /w:[ 1 0 7 0 ]
  //: joint g17 (Reset) @(467, 308) /w:[ 5 -1 6 8 ]
  _GGNAND2 #(4) g2 (.I0(w2), .I1(w7), .Z(w8));   //: @(402,212) /sn:0 /w:[ 1 5 5 ]
  //: joint g23 (Q) @(650, 218) /w:[ 5 -1 6 8 ]
  //: joint g24 (Qinv) @(670, 270) /w:[ 1 2 4 -1 ]
  _GGNAND3 #(6) g1 (.I0(CLK), .I1(Q), .I2(K), .Z(w5));   //: @(310,274) /sn:0 /w:[ 9 0 1 0 ]
  //: joint g18 (Reset) @(589, 308) /w:[ -1 2 4 1 ]
  //: joint g25 (Q) @(682, 218) /w:[ 2 -1 4 1 ]
  //: IN g10 (K) @(178,279) /sn:0 /w:[ 0 ]
  _GGNAND2 #(4) g6 (.I0(w14), .I1(Qinv), .Z(Q));   //: @(619,218) /sn:0 /w:[ 1 7 7 ]
  _GGNAND3 #(6) g7 (.I0(Q), .I1(w13), .I2(Reset), .Z(Qinv));   //: @(619,270) /sn:0 /w:[ 9 1 3 9 ]
  //: IN g9 (J) @(183,205) /sn:0 /w:[ 0 ]
  //: joint g22 (Qinv) @(659, 270) /w:[ 5 6 8 -1 ]
  //: IN g12 (Reset) @(467,360) /sn:0 /R:1 /w:[ 9 ]
  _GGNAND2 #(4) g5 (.I0(w26), .I1(w7), .Z(w13));   //: @(524,270) /sn:0 /w:[ 3 3 0 ]
  //: OUT g14 (Qinv) @(707,270) /sn:0 /w:[ 0 ]
  //: IN g11 (CLK) @(195,335) /sn:0 /w:[ 0 ]
  //: joint g21 (w8) @(434, 212) /w:[ 2 -1 4 1 ]
  //: joint g19 (w26) @(488, 267) /w:[ 2 1 -1 4 ]
  //: joint g20 (w7) @(450, 279) /w:[ 2 4 1 -1 ]
  _GGNAND3 #(6) g0 (.I0(J), .I1(Qinv), .I2(CLK), .Z(w2));   //: @(312,210) /sn:0 /w:[ 1 3 11 0 ]
  //: joint g15 (CLK) @(293, 335) /w:[ 2 4 1 6 ]
  //: OUT g13 (Q) @(703,217) /sn:0 /w:[ 3 ]

endmodule
//: /netlistEnd

