//: version "2.1"
//: property encoding = "utf-8"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "Lab5_A.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg CLOCK;    //: /sn:0 {0}(338,232)(320,232){1}
//: {2}(316,232)(272,232){3}
//: {4}(268,232)(246,232){5}
//: {6}(244,230)(244,65)(308,65){7}
//: {8}(310,63)(310,3)(343,3){9}
//: {10}(310,67)(310,126)(341,126){11}
//: {12}(242,232)(155,232){13}
//: {14}(151,232)(13:83,232){15}
//: {16}(153,234)(153,428)(316,428){17}
//: {18}(270,234)(270,277){19}
//: {20}(318,234)(318,237)(338,237){21}
reg K;    //: /sn:0 {0}(97:341,131)(124,131){1}
//: {2}(120,131)(81,131){3}
//: {4}(122,133)(122,462)(316,462){5}
reg J;    //: /sn:0 {0}(80:79,-2)(197,-2){1}
//: {2}(201,-2)(343,-2){3}
//: {4}(199,0)(199,396)(316,396){5}
reg Reset;    //: /sn:0 {0}(383,496)(383,558)(583,558)(583,301)(384,301){1}
//: {2}(382,299)(382,166){3}
//: {4}(384,164)(562,164)(562,134)(577,134){5}
//: {6}(382,162)(382,136)(399,136){7}
//: {8}(382,303)(1:382,316){9}
wire w6;    //: /sn:0 {0}(399,131)(362,131){1}
wire w13;    //: /sn:0 {0}(453,447)(485,447)(485,426){1}
wire w7;    //: /sn:0 {0}(594,5)(613,5){1}
//: {2}(617,5)(654,5){3}
//: {4}(658,5)(726,5)(726,-9){5}
//: {6}(656,7)(656,184)(324,184)(324,136)(341,136){7}
//: {8}(615,7)(615,86)(566,86)(566,124)(577,124){9}
wire w4;    //: /sn:0 {0}(429,-54)(429,-3){1}
//: {2}(431,-1)(521,-1){3}
//: {4}(427,-1)(402,-1){5}
//: {6}(429,1)(429,100)(382,100)(382,126)(399,126){7}
wire w0;    //: /sn:0 {0}(573,7)(563,7)(563,64)(629,64)(629,127){1}
//: {2}(631,129)(685,129)(685,-21)(328,-21)(328,-7)(343,-7){3}
//: {4}(627,129)(598,129){5}
wire w10;    //: /sn:0 {0}(577,129)(540,129){1}
wire w1;    //: /sn:0 {0}(454,268)(454,237){1}
//: {2}(456,235)(474,235)(474,69)(502,69){3}
//: {4}(504,67)(504,4)(521,4){5}
//: {6}(504,71)(504,126)(519,126){7}
//: {8}(452,235)(359,235){9}
wire w8;    //: /sn:0 {0}(573,2)(542,2){1}
wire w14;    //: /sn:0 {0}(453,406)(468,406)(468,382){1}
wire w2;    //: /sn:0 {0}(381,-3)(366,-3)(366,-2)(364,-2){1}
wire w5;    //: /sn:0 {0}(519,131)(450,131){1}
//: {2}(448,129)(448,61)(377,61)(377,2)(381,2){3}
//: {4}(446,131)(420,131){5}
//: enddecls

  _GGNAND2 #(4) g4 (.I0(w2), .I1(w5), .Z(w4));   //: @(392,-1) /sn:0 /w:[ 0 3 5 ]
  //: joint g8 (CLOCK) @(244, 232) /w:[ 5 6 12 -1 ]
  //: joint g16 (w7) @(615, 5) /w:[ 2 -1 1 8 ]
  _GGNAND3 #(6) g3 (.I0(CLOCK), .I1(K), .I2(w7), .Z(w6));   //: @(352,131) /sn:0 /w:[ 11 0 7 1 ]
  //: LED Qs (w7) @(726,-16) /sn:0 /w:[ 5 ] /type:0
  //: joint g17 (CLOCK) @(270, 232) /w:[ 3 -1 4 18 ]
  //: comment g26 @(368,346) /sn:0
  //: /line:"RESET"
  //: /end
  //: LED Qm (w4) @(429,-61) /sn:0 /w:[ 0 ] /type:0
  _GGNAND3 #(6) g2 (.I0(w0), .I1(J), .I2(CLOCK), .Z(w2));   //: @(354,-2) /sn:0 /w:[ 3 3 9 1 ]
  //: joint g23 (w1) @(454, 235) /w:[ 2 -1 8 1 ]
  //: comment g30 @(736,-24) /sn:0
  //: /line:"Qs"
  //: /end
  //: SWITCH g1 (K) @(64,131) /sn:0 /w:[ 3 ] /st:0 /dn:0
  //: LED g24 (w1) @(454,275) /sn:0 /R:2 /w:[ 0 ] /type:0
  //: comment g29 @(89,214) /sn:0
  //: /line:"CLOCK"
  //: /end
  _GGNAND2 #(4) g18 (.I0(CLOCK), .I1(CLOCK), .Z(w1));   //: @(349,235) /sn:0 /w:[ 0 21 9 ]
  _GGNAND2 #(4) g10 (.I0(w1), .I1(w5), .Z(w10));   //: @(530,129) /sn:0 /w:[ 7 0 1 ]
  //: SWITCH J1 (J) @(62,-3) /sn:0 /w:[ 0 ] /st:0 /dn:0
  //: joint g25 (Reset) @(382, 164) /w:[ 4 6 -1 3 ]
  //: joint g6 (w4) @(429, -1) /w:[ 2 1 4 6 ]
  //: LED g35 (w13) @(485,419) /sn:0 /w:[ 1 ] /type:0
  _GGNAND2 #(4) g9 (.I0(w4), .I1(w1), .Z(w8));   //: @(532,2) /sn:0 /w:[ 3 5 1 ]
  //: joint g7 (w5) @(448, 131) /w:[ 1 2 4 -1 ]
  //: SWITCH g22 (Reset) @(382,330) /sn:0 /R:1 /w:[ 9 ] /st:1 /dn:0
  //: comment g31 @(439,-66) /sn:0
  //: /line:"Qm"
  //: /end
  //: joint g33 (Reset) @(382, 301) /w:[ 1 2 -1 8 ]
  //: joint g36 (J) @(199, -2) /w:[ 2 -1 1 4 ]
  _GGNAND3 #(6) g12 (.I0(w7), .I1(w10), .I2(Reset), .Z(w0));   //: @(588,129) /sn:0 /w:[ 9 0 5 5 ]
  //: LED g34 (w14) @(468,375) /sn:0 /w:[ 1 ] /type:0
  //: comment g28 @(89,112) /sn:0
  //: /line:"K"
  //: /end
  _GGNAND2 #(4) g11 (.I0(w8), .I1(w0), .Z(w7));   //: @(584,5) /sn:0 /w:[ 0 0 0 ]
  _GGNAND3 #(6) g5 (.I0(w4), .I1(w6), .I2(Reset), .Z(w5));   //: @(410,131) /sn:0 /w:[ 7 0 7 5 ]
  //: joint g14 (CLOCK) @(310, 65) /w:[ -1 8 7 10 ]
  //: LED g19 (CLOCK) @(270,284) /sn:0 /R:2 /w:[ 19 ] /type:0
  //: joint g21 (w1) @(504, 69) /w:[ -1 4 3 6 ]
  //: joint g20 (CLOCK) @(318, 232) /w:[ 1 -1 2 20 ]
  JKFlipFlop g32 (.J(J), .K(K), .CLOCK(CLOCK), .RESET(Reset), .Q(w14), .Qinv(w13));   //: @(317, 377) /sz:(135, 118) /sn:0 /p:[ Li0>5 Li1>5 Li2>17 Bi0>0 Ro0<0 Ro1<0 ]
  //: joint g15 (w0) @(629, 129) /w:[ 2 1 4 -1 ]
  //: SWITCH g0 (CLOCK) @(66,232) /sn:0 /w:[ 15 ] /st:0 /dn:0
  //: joint g38 (CLOCK) @(153, 232) /w:[ 13 -1 14 16 ]
  //: comment g27 @(87,-20) /sn:0
  //: /line:"<big>J</big>"
  //: /end
  //: joint g37 (K) @(122, 131) /w:[ 1 -1 2 4 ]
  //: joint g13 (w7) @(656, 5) /w:[ 4 -1 3 6 ]

endmodule
//: /netlistEnd

//: /netlistBegin JKFlipFlop
module JKFlipFlop(CLOCK, RESET, K, Q, Qinv, J);
//: interface  /sz:(135, 118) /bd:[ Li0>J(19/118) Li1>K(85/118) Li2>CLOCK(51/118) Bi0>RESET(66/135) Ro0<Q(29/118) Ro1<Qinv(70/118) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input CLOCK;    //: /sn:0 {0}(256,222)(240,222)(240,253){1}
//: {2}(238,255)(227,255)(227,348){3}
//: {4}(229,350)(242,350){5}
//: {6}(246,350)(256,350){7}
//: {8}(244,352)(244,355)(256,355){9}
//: {10}(225,350)(205,350){11}
//: {12}(240,257)(240,288)(255,288){13}
output Q;    //: /sn:0 {0}(642,226)(578,226)(578,226)(602,226){1}
//: {2}(598,226)(542,226){3}
//: {4}(538,226)(524,226){5}
//: {6}(540,228)(540,258)(486,258)(486,286)(506,286){7}
//: {8}(600,228)(600,330)(242,330)(242,298)(255,298){9}
input K;    //: /sn:0 {0}(255,293)(239,293)(239,293)(204,293){1}
input RESET;    //: /sn:0 {0}(382,380)(382,321){1}
//: {2}(384,319)(491,319)(491,296)(506,296){3}
//: {4}(380,319)(331,319)(331,298)(346,298){5}
output Qinv;    //: /sn:0 {0}(640,291)(609,291)(609,291)(588,291){1}
//: {2}(586,289)(586,177)(230,177)(230,212)(256,212){3}
//: {4}(584,291)(571,291){5}
//: {6}(569,289)(569,251)(494,251)(494,228)(503,228){7}
//: {8}(567,291)(564,291)(564,291)(527,291){9}
input J;    //: /sn:0 {0}(256,217)(241,217)(241,217)(208,217){1}
wire w6;    //: /sn:0 {0}(346,293)(330,293)(330,293)(276,293){1}
wire w7;    //: /sn:0 {0}(458,293)(443,293)(443,293)(393,293){1}
//: {2}(391,291)(391,255)(328,255)(328,222)(352,222){3}
//: {4}(389,293)(367,293){5}
wire w4;    //: /sn:0 {0}(451,220)(430,220)(430,220)(387,220){1}
//: {2}(383,220)(373,220){3}
//: {4}(385,222)(385,262)(319,262)(319,288)(346,288){5}
wire w14;    //: /sn:0 {0}(479,291)(494,291)(494,291)(506,291){1}
wire w2;    //: /sn:0 {0}(352,217)(303,217)(303,217)(277,217){1}
wire w5;    //: /sn:0 {0}(503,223)(488,223)(488,223)(472,223){1}
wire w9;    //: /sn:0 {0}(458,288)(438,288)(438,257){1}
//: {2}(438,253)(438,225)(451,225){3}
//: {4}(436,255)(420,255)(420,353)(277,353){5}
//: enddecls

  _GGNAND3 #(6) g4 (.I0(CLOCK), .I1(K), .I2(Q), .Z(w6));   //: @(266,293) /sn:0 /w:[ 13 0 9 1 ]
  //: joint g8 (CLOCK) @(244, 350) /w:[ 6 -1 5 8 ]
  _GGNAND3 #(6) g3 (.I0(Qinv), .I1(J), .I2(CLOCK), .Z(w2));   //: @(267,217) /sn:0 /w:[ 3 0 0 1 ]
  _GGNAND3 #(6) g16 (.I0(Q), .I1(w14), .I2(RESET), .Z(Qinv));   //: @(517,291) /sn:0 /w:[ 7 1 3 9 ]
  //: joint g17 (Q) @(540, 226) /w:[ 3 -1 4 6 ]
  //: IN g2 (CLOCK) @(203,350) /sn:0 /w:[ 11 ]
  //: IN g23 (RESET) @(382,382) /sn:0 /R:1 /w:[ 0 ]
  //: IN g1 (K) @(202,293) /sn:0 /w:[ 1 ]
  //: OUT g24 (Q) @(639,226) /sn:0 /w:[ 0 ]
  //: joint g18 (Qinv) @(569, 291) /w:[ 5 6 8 -1 ]
  //: joint g10 (CLOCK) @(227, 350) /w:[ 4 3 10 -1 ]
  //: OUT g25 (Qinv) @(637,291) /sn:0 /w:[ 0 ]
  _GGNAND2 #(4) g6 (.I0(w2), .I1(w7), .Z(w4));   //: @(363,220) /sn:0 /w:[ 0 3 3 ]
  _GGNAND3 #(6) g7 (.I0(w4), .I1(w6), .I2(RESET), .Z(w7));   //: @(357,293) /sn:0 /w:[ 5 0 5 5 ]
  //: joint g9 (CLOCK) @(240, 255) /w:[ -1 1 2 12 ]
  //: joint g22 (Q) @(600, 226) /w:[ 1 -1 2 8 ]
  //: joint g12 (w4) @(385, 220) /w:[ 1 -1 2 4 ]
  _GGNAND2 #(4) g5 (.I0(CLOCK), .I1(CLOCK), .Z(w9));   //: @(267,353) /sn:0 /w:[ 7 9 5 ]
  //: joint g11 (w7) @(391, 293) /w:[ 1 2 4 -1 ]
  _GGNAND2 #(4) g14 (.I0(w5), .I1(Qinv), .Z(Q));   //: @(514,226) /sn:0 /w:[ 0 7 5 ]
  //: joint g21 (Qinv) @(586, 291) /w:[ 1 2 4 -1 ]
  //: joint g19 (RESET) @(382, 319) /w:[ 2 -1 4 1 ]
  //: joint g20 (w9) @(438, 255) /w:[ -1 2 4 1 ]
  //: IN g0 (J) @(206,217) /sn:0 /w:[ 1 ]
  _GGNAND2 #(4) g15 (.I0(w9), .I1(w7), .Z(w14));   //: @(469,291) /sn:0 /w:[ 0 0 0 ]
  _GGNAND2 #(4) g13 (.I0(w4), .I1(w9), .Z(w5));   //: @(462,223) /sn:0 /w:[ 0 3 1 ]

endmodule
//: /netlistEnd

