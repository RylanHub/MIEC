//: version "2.1"
//: property encoding = "utf-8"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "Lab4_B.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
supply1 w6;    //: /sn:0 {0}(628,343)(346,343)(346,318){1}
//: {2}(348,316)(628,316){3}
//: {4}(346,314)(346,132){5}
reg B;    //: /sn:0 {0}(522,593)(522,496){1}
supply0 w4;    //: /sn:0 {0}(324,439)(324,325){1}
//: {2}(326,323)(628,323){3}
//: {4}(324,321)(324,305){5}
//: {6}(326,303)(628,303){7}
//: {8}(324,301)(324,296)(628,296){9}
reg A;    //: /sn:0 {0}(357,565)(357,558)(512,558)(512,496){1}
reg D;    //: /sn:0 {0}(204,310)(217,310){1}
//: {2}(221,310)(234,310){3}
//: {4}(238,310)(628,310){5}
//: {6}(236,312)(236,336)(628,336){7}
//: {8}(219,312)(219,330)(628,330){9}
reg C;    //: /sn:0 {0}(532,496)(532,557)(592,557)(592,570){1}
wire [2:0] w15;    //: /sn:0 {0}(644,343)(644,418)(522,418)(#:522,490){1}
wire w9;    //: /sn:0 {0}(657,320)(691,320)(691,279){1}
//: enddecls

  //: VDD g8 (w6) @(357,132) /sn:0 /w:[ 5 ]
  //: SWITCH g4 (C) @(592,584) /sn:0 /R:1 /w:[ 1 ] /st:1 /dn:1
  //: SWITCH g3 (B) @(522,607) /sn:0 /R:1 /w:[ 0 ] /st:0 /dn:1
  _GGMUX8 #(20, 22) g2 (.I0(w6), .I1(D), .I2(D), .I3(w4), .I4(w6), .I5(~D), .I6(w4), .I7(w4), .S(w15), .Z(w9));   //: @(644,320) /sn:0 /R:1 /w:[ 0 7 9 3 3 5 7 9 0 0 ] /ss:0 /do:0
  //: SWITCH g1 (A) @(357,579) /sn:0 /R:1 /w:[ 0 ] /st:1 /dn:1
  //: joint g10 (D) @(219, 310) /w:[ 2 -1 1 8 ]
  //: GROUND g6 (w4) @(324,445) /sn:0 /w:[ 0 ]
  //: joint g9 (w6) @(346, 316) /w:[ 2 4 -1 1 ]
  //: SWITCH g7 (D) @(187,310) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: LED g12 (w9) @(691,272) /sn:0 /w:[ 1 ] /type:0
  //: joint g11 (D) @(236, 310) /w:[ 4 -1 3 6 ]
  //: joint g5 (w4) @(324, 303) /w:[ 6 8 -1 5 ]
  assign w15 = {A, B, C}; //: CONCAT g0  @(522,491) /sn:0 /R:1 /w:[ 1 1 1 0 ] /dr:0 /tp:0 /drp:1
  //: joint g13 (w4) @(324, 323) /w:[ 2 4 -1 1 ]

endmodule
//: /netlistEnd

