//: version "2.1"
//: property encoding = "utf-8"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "Lab3_A.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg B;    //: /sn:0 {0}(584,244)(581,244)(581,296)(521,296){1}
//: {2}(517,296)(458,296){3}
//: {4}(454,296)(328,296){5}
//: {6}(456,298)(456,348)(585,348){7}
//: {8}(519,298)(519,417)(588,417){9}
reg A;    //: /sn:0 {0}(584,239)(568,239)(568,220)(497,220){1}
//: {2}(493,220)(402,220){3}
//: {4}(398,220)(329,220){5}
//: {6}(400,222)(400,343)(585,343){7}
//: {8}(495,222)(495,412)(588,412){9}
reg D;    //: /sn:0 {0}(586,461)(448,461){1}
//: {2}(446,459)(446,353)(585,353){3}
//: {4}(444,461)(334,461){5}
reg C;    //: /sn:0 {0}(588,422)(468,422)(468,379){1}
//: {2}(470,377)(579,377)(579,456)(586,456){3}
//: {4}(466,377)(388,377){5}
//: {6}(386,375)(386,249)(584,249){7}
//: {8}(384,377)(334,377){9}
wire w6;    //: /sn:0 {0}(607,459)(680,459)(680,358)(693,358){1}
wire w4;    //: /sn:0 {0}(693,353)(678,353)(678,417)(609,417){1}
wire w3;    //: /sn:0 {0}(693,348)(606,348){1}
wire w2;    //: /sn:0 {0}(693,343)(678,343)(678,244)(605,244){1}
wire w5;    //: /sn:0 {0}(728,335)(728,350)(714,350){1}
//: enddecls

  //: joint g8 (A) @(400, 220) /w:[ 3 -1 4 6 ]
  _GGAND3 #(8) g4 (.I0(!A), .I1(B), .I2(!C), .Z(w2));   //: @(595,244) /sn:0 /w:[ 0 0 7 1 ]
  //: LED g16 (w5) @(728,328) /sn:0 /w:[ 0 ] /type:0
  //: SWITCH g3 (D) @(317,461) /sn:0 /w:[ 5 ] /st:1 /dn:1
  //: SWITCH g2 (C) @(317,377) /sn:0 /w:[ 9 ] /st:0 /dn:1
  //: SWITCH g1 (B) @(311,296) /sn:0 /w:[ 5 ] /st:1 /dn:1
  //: joint g10 (D) @(446, 461) /w:[ 1 2 4 -1 ]
  //: joint g6 (C) @(386, 377) /w:[ 5 6 8 -1 ]
  //: joint g9 (B) @(456, 296) /w:[ 3 -1 4 6 ]
  _GGAND3 #(8) g7 (.I0(A), .I1(!B), .I2(!D), .Z(w3));   //: @(596,348) /sn:0 /w:[ 7 7 3 1 ]
  //: joint g12 (A) @(495, 220) /w:[ 1 -1 2 8 ]
  //: joint g14 (C) @(468, 377) /w:[ 2 -1 4 1 ]
  _GGAND3 #(8) g11 (.I0(A), .I1(!B), .I2(!C), .Z(w4));   //: @(599,417) /sn:0 /w:[ 9 9 0 1 ]
  _GGAND2 #(4) g5 (.I0(!C), .I1(!D), .Z(w6));   //: @(597,459) /sn:0 /w:[ 3 0 0 ]
  _GGOR4 #(10) g15 (.I0(w2), .I1(w3), .I2(w4), .I3(w6), .Z(w5));   //: @(704,350) /sn:0 /w:[ 0 0 0 1 1 ]
  //: SWITCH g0 (A) @(312,220) /sn:0 /w:[ 5 ] /st:0 /dn:1
  //: joint g13 (B) @(519, 296) /w:[ 1 -1 2 8 ]

endmodule
//: /netlistEnd

