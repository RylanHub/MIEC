//: version "2.1"
//: property encoding = "utf-8"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "Lab5_A.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg CLOCK;    //: /sn:0 {0}(301,397)(283,397){1}
//: {2}(279,397)(235,397){3}
//: {4}(231,397)(209,397){5}
//: {6}(207,395)(207,230)(271,230){7}
//: {8}(273,228)(273,168)(306,168){9}
//: {10}(273,232)(273,291)(304,291){11}
//: {12}(205,397)(13:137,397){13}
//: {14}(233,399)(233,442){15}
//: {16}(281,399)(281,402)(301,402){17}
reg K;    //: /sn:0 {0}(97:304,296)(136,296){1}
reg J;    //: /sn:0 {0}(306,163)(80:133,163){1}
reg Reset;    //: /sn:0 {0}(1:345,430)(345,331){1}
//: {2}(347,329)(525,329)(525,299)(540,299){3}
//: {4}(345,327)(345,301)(362,301){5}
wire w6;    //: /sn:0 {0}(362,296)(325,296){1}
wire w7;    //: /sn:0 {0}(557,171)(577,171){1}
//: {2}(581,171)(619,171){3}
//: {4}(623,171)(689,171)(689,156){5}
//: {6}(621,173)(621,350)(289,350)(289,301)(304,301){7}
//: {8}(579,173)(579,252)(530,252)(530,289)(540,289){9}
wire w4;    //: /sn:0 {0}(484,165)(396,165){1}
//: {2}(394,163)(394,116){3}
//: {4}(392,165)(378,165){5}
//: {6}(394,167)(394,256)(343,256)(343,291)(362,291){7}
wire w0;    //: /sn:0 {0}(536,173)(526,173)(526,230)(592,230)(592,292){1}
//: {2}(594,294)(648,294)(648,144)(291,144)(291,158)(306,158){3}
//: {4}(590,294)(561,294){5}
wire w10;    //: /sn:0 {0}(540,294)(503,294){1}
wire w1;    //: /sn:0 {0}(417,433)(417,402){1}
//: {2}(419,400)(437,400)(437,234)(465,234){3}
//: {4}(467,232)(467,170)(484,170){5}
//: {6}(467,236)(467,291)(482,291){7}
//: {8}(415,400)(322,400){9}
wire w8;    //: /sn:0 {0}(536,168)(505,168){1}
wire w2;    //: /sn:0 {0}(357,163)(327,163){1}
wire w5;    //: /sn:0 {0}(482,296)(413,296){1}
//: {2}(411,294)(411,227)(353,227)(353,168)(357,168){3}
//: {4}(409,296)(383,296){5}
//: enddecls

  //: joint g8 (CLOCK) @(207, 397) /w:[ 5 6 12 -1 ]
  _GGNAND2 #(4) g4 (.I0(w2), .I1(w5), .Z(w4));   //: @(368,165) /sn:0 /w:[ 0 3 5 ]
  _GGNAND3 #(6) g3 (.I0(CLOCK), .I1(K), .I2(w7), .Z(w6));   //: @(315,296) /sn:0 /w:[ 11 0 7 1 ]
  //: joint g16 (w7) @(579, 171) /w:[ 2 -1 1 8 ]
  //: comment g26 @(331,460) /sn:0
  //: /line:"RESET"
  //: /end
  //: joint g17 (CLOCK) @(233, 397) /w:[ 3 -1 4 14 ]
  //: LED Qs (w7) @(689,149) /sn:0 /w:[ 5 ] /type:0
  _GGNAND3 #(6) g2 (.I0(w0), .I1(J), .I2(CLOCK), .Z(w2));   //: @(317,163) /sn:0 /w:[ 3 0 9 1 ]
  //: LED Qm (w4) @(394,109) /sn:0 /w:[ 3 ] /type:0
  //: comment g30 @(699,141) /sn:0
  //: /line:"Qs"
  //: /end
  //: joint g23 (w1) @(417, 400) /w:[ 2 -1 8 1 ]
  //: LED g24 (w1) @(417,440) /sn:0 /R:2 /w:[ 0 ] /type:0
  //: SWITCH g1 (K) @(119,296) /sn:0 /w:[ 1 ] /st:1 /dn:0
  //: comment g29 @(143,379) /sn:0
  //: /line:"CLOCK"
  //: /end
  _GGNAND2 #(4) g18 (.I0(CLOCK), .I1(CLOCK), .Z(w1));   //: @(312,400) /sn:0 /w:[ 0 17 9 ]
  //: joint g25 (Reset) @(345, 329) /w:[ 2 4 -1 1 ]
  //: SWITCH J1 (J) @(116,162) /sn:0 /w:[ 1 ] /st:0 /dn:0
  _GGNAND2 #(4) g10 (.I0(w1), .I1(w5), .Z(w10));   //: @(493,294) /sn:0 /w:[ 7 0 1 ]
  //: joint g6 (w4) @(394, 165) /w:[ 1 2 4 6 ]
  //: joint g7 (w5) @(411, 296) /w:[ 1 2 4 -1 ]
  _GGNAND2 #(4) g9 (.I0(w4), .I1(w1), .Z(w8));   //: @(495,168) /sn:0 /w:[ 0 5 1 ]
  //: comment g31 @(404,101) /sn:0
  //: /line:"Qm"
  //: /end
  //: SWITCH g22 (Reset) @(345,444) /sn:0 /R:1 /w:[ 0 ] /st:1 /dn:0
  _GGNAND3 #(6) g12 (.I0(w7), .I1(w10), .I2(Reset), .Z(w0));   //: @(551,294) /sn:0 /w:[ 9 0 3 5 ]
  //: comment g28 @(143,277) /sn:0
  //: /line:"K"
  //: /end
  //: joint g14 (CLOCK) @(273, 230) /w:[ -1 8 7 10 ]
  _GGNAND3 #(6) g5 (.I0(w4), .I1(w6), .I2(Reset), .Z(w5));   //: @(373,296) /sn:0 /w:[ 7 0 5 5 ]
  _GGNAND2 #(4) g11 (.I0(w8), .I1(w0), .Z(w7));   //: @(547,171) /sn:0 /w:[ 0 0 0 ]
  //: joint g21 (w1) @(467, 234) /w:[ -1 4 3 6 ]
  //: LED g19 (CLOCK) @(233,449) /sn:0 /R:2 /w:[ 15 ] /type:0
  //: joint g20 (CLOCK) @(281, 397) /w:[ 1 -1 2 16 ]
  //: SWITCH g0 (CLOCK) @(120,397) /sn:0 /w:[ 13 ] /st:0 /dn:0
  //: joint g15 (w0) @(592, 294) /w:[ 2 1 4 -1 ]
  //: comment g27 @(141,145) /sn:0
  //: /line:"<big>J</big>"
  //: /end
  //: joint g13 (w7) @(621, 171) /w:[ 4 -1 3 6 ]

endmodule
//: /netlistEnd

//: /netlistBegin JKFlipFlop
module JKFlipFlop();
//: interface  /sz:(135, 118) /bd:[ Li0>CLOCK(51/118) Li1>K(85/118) Li2>J(19/118) Bi0>RESET(66/135) Ro0<Qinv(70/118) Ro1<Q(29/118) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
//: enddecls


endmodule
//: /netlistEnd

