//: version "2.1"
//: property encoding = "utf-8"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "Lab3.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg X;    //: /sn:0 {0}(112,88)(139,88){1}
//: {2}(143,88)(183,88)(183,115)(196,115){3}
//: {4}(141,90)(141,208)(199,208){5}
reg Z;    //: /sn:0 {0}(114,248)(309,248)(309,196){1}
//: {2}(311,194)(438,194){3}
//: {4}(309,192)(309,152)(440,152){5}
reg Y;    //: /sn:0 {0}(196,120)(181,120)(181,136)(129,136){1}
//: {2}(125,136)(115,136){3}
//: {4}(127,138)(127,213)(199,213){5}
wire w3;    //: /sn:0 {0}(475,134)(475,150)(461,150){1}
wire w12;    //: /sn:0 {0}(523,179)(523,209)(522,209){1}
wire w2;    //: /sn:0 {0}(440,147)(409,147)(409,118)(376,118){1}
//: {2}(372,118)(217,118){3}
//: {4}(374,120)(374,189)(438,189){5}
wire w5;    //: /sn:0 {0}(220,211)(501,211){1}
wire w9;    //: /sn:0 {0}(501,206)(487,206)(487,192)(459,192){1}
//: enddecls

  //: joint g4 (X) @(141, 88) /w:[ 2 -1 1 4 ]
  _GGAND2 #(6) g8 (.I0(w2), .I1(Z), .Z(w9));   //: @(449,192) /sn:0 /w:[ 5 3 1 ]
  //: SWITCH X (X) @(95,88) /sn:0 /w:[ 0 ] /st:1 /dn:1
  //: joint g2 (Y) @(127, 136) /w:[ 1 -1 2 4 ]
  _GGAND2 #(6) g1 (.I0(X), .I1(Y), .Z(w5));   //: @(210,211) /sn:0 /w:[ 5 5 0 ]
  //: LED carry (w12) @(523,172) /w:[ 0 ] /type:0
  //: joint g10 (w2) @(374, 118) /w:[ 1 -1 2 4 ]
  _GGXOR2 #(8) g6 (.I0(w2), .I1(Z), .Z(w3));   //: @(451,150) /sn:0 /w:[ 0 5 1 ]
  //: SWITCH g7 (Z) @(97,248) /sn:0 /w:[ 0 ] /st:0 /dn:1
  _GGOR2 #(6) g9 (.I0(w9), .I1(w5), .Z(w12));   //: @(512,209) /sn:0 /w:[ 0 1 1 ]
  //: joint g11 (Z) @(309, 194) /w:[ 2 4 -1 1 ]
  //: LED sum (w3) @(475,127) /w:[ 0 ] /type:0
  _GGXOR2 #(8) g0 (.I0(X), .I1(Y), .Z(w2));   //: @(207,118) /sn:0 /w:[ 3 0 3 ]
  //: SWITCH Y (Y) @(98,136) /sn:0 /w:[ 3 ] /st:1 /dn:1

endmodule
//: /netlistEnd

