//: version "2.1"
//: property encoding = "utf-8"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "Lab6.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg [3:0] B;    //: /sn:0 {0}(#:268,291)(204,291)(#:204,271){1}
reg [3:0] A;    //: /sn:0 {0}(#:274,135)(208,135)(#:208,114){1}
supply0 w17;    //: /sn:0 {0}(426,89)(426,35){1}
wire w13;    //: /sn:0 {0}(663,258)(710,258)(710,237)(783,237){1}
wire w6;    //: /sn:0 {0}(274,278)(345,278)(345,258)(385,258){1}
wire w7;    //: /sn:0 {0}(385,282)(347,282)(347,288)(274,288){1}
wire w4;    //: /sn:0 {0}(385,145)(355,145)(355,142)(280,142){1}
wire w3;    //: /sn:0 {0}(385,127)(355,127)(355,132)(280,132){1}
wire w12;    //: /sn:0 {0}(663,227)(783,227){1}
wire w10;    //: /sn:0 {0}(663,164)(714,164)(714,207)(725,207)(783,207){1}
wire w8;    //: /sn:0 {0}(385,305)(348,305)(348,298)(274,298){1}
wire w14;    //: /sn:0 {0}(663,287)(716,287)(716,247)(783,247){1}
wire w11;    //: /sn:0 {0}(783,217)(703,217)(703,193)(663,193){1}
wire w2;    //: /sn:0 {0}(280,122)(355,122)(355,108)(385,108){1}
wire [4:0] w15;    //: /sn:0 {0}(818,145)(818,227)(#:789,227){1}
wire w5;    //: /sn:0 {0}(385,164)(354,164)(354,152)(280,152){1}
wire w9;    //: /sn:0 {0}(385,327)(344,327)(344,308)(274,308){1}
//: enddecls

  assign {w9, w8, w7, w6} = B; //: CONCAT g4  @(269,293) /sn:0 /R:2 /w:[ 1 1 1 0 0 ] /dr:0 /tp:0 /drp:0
  //: comment g8 @(150,183) /sn:0
  //: /line:"4-bit number A and B"
  //: /line:"ranging from 0 to F "
  //: /line:"in hexadecimal form"
  //: /end
  //: GROUND g3 (w17) @(426,29) /sn:0 /R:2 /w:[ 1 ]
  assign {w5, w4, w3, w2} = A; //: CONCAT g2  @(275,137) /sn:0 /R:2 /w:[ 1 1 1 0 0 ] /dr:0 /tp:0 /drp:0
  LookAheadAdder g1 (.cin(w17), .a0(w2), .a1(w3), .a2(w4), .a3(w5), .b0(w6), .b1(w7), .b2(w8), .b3(w9), .cout(w14), .s0(w10), .s1(w11), .s2(w12), .s3(w13));   //: @(386, 90) /sz:(276, 260) /sn:0 /p:[ Ti0>0 Li0>1 Li1>0 Li2>0 Li3>0 Li4>1 Li5>0 Li6>0 Li7>0 Ro0<0 Ro1<0 Ro2<1 Ro3<0 Ro4<0 ]
  assign w15 = {w14, w13, w12, w11, w10}; //: CONCAT g6  @(788,227) /sn:0 /w:[ 1 1 1 1 0 1 ] /dr:1 /tp:0 /drp:1
  //: LED g7 (w15) @(818,138) /sn:0 /w:[ 0 ] /type:3
  //: comment g9 @(761,59) /sn:0
  //: /line:"5-bit sum"
  //: /line:"ranging from 0 to 31 "
  //: /line:"in decimal form"
  //: /end
  //: DIP g5 (B) @(204,261) /sn:0 /w:[ 1 ] /st:14 /dn:1
  //: DIP g0 (A) @(208,104) /sn:0 /w:[ 1 ] /st:13 /dn:1

endmodule
//: /netlistEnd

//: /netlistBegin LookAheadAdder
module LookAheadAdder(b0, cin, a0, cout, a2, b3, a3, b1, s1, s2, a1, s0, b2, s3);
//: interface  /sz:(276, 260) /bd:[ Ti0>cin(40/276) Li0>a0(18/260) Li1>a1(37/260) Li2>a2(55/260) Li3>a3(74/260) Li4>b0(168/260) Li5>b1(192/260) Li6>b2(215/260) Li7>b3(237/260) Ro0<cout(197/260) Ro1<s0(74/260) Ro2<s1(103/260) Ro3<s2(137/260) Ro4<s3(168/260) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output s2;    //: /sn:0 {0}(-16,376)(-16,366)(-16,366)(-16,367){1}
input a2;    //: /sn:0 {0}(-16,346)(-16,156){1}
//: {2}(-14,154)(122,154){3}
//: {4}(126,154)(142,154){5}
//: {6}(124,156)(124,211)(139,211){7}
//: {8}(-18,154)(-126,154){9}
output s0;    //: /sn:0 {0}(-106,376)(-106,365)(-106,365)(-106,365){1}
input b2;    //: /sn:0 {0}(-126,159)(-13,159){1}
//: {2}(-9,159)(107,159){3}
//: {4}(111,159)(142,159){5}
//: {6}(109,161)(109,216)(139,216){7}
//: {8}(-11,161)(-11,346){9}
input a3;    //: /sn:0 {0}(-127,256)(-39,256)(-39,256)(33,256){1}
//: {2}(37,256)(86,256)(86,256)(121,256){3}
//: {4}(125,256)(141,256){5}
//: {6}(123,258)(123,341)(139,341){7}
//: {8}(35,258)(35,345){9}
input b3;    //: /sn:0 {0}(-127,261)(38,261){1}
//: {2}(42,261)(106,261){3}
//: {4}(110,261)(141,261){5}
//: {6}(108,263)(108,346)(139,346){7}
//: {8}(40,263)(40,345){9}
output s3;    //: /sn:0 {0}(35,376)(35,366)(35,366)(35,366){1}
output s1;    //: /sn:0 {0}(-60,366)(-60,366)(-60,366)(-60,376){1}
input a1;    //: /sn:0 {0}(141,76)(133,76)(133,76)(129,76){1}
//: {2}(125,76)(-58,76){3}
//: {4}(-62,76)(-123,76){5}
//: {6}(-60,78)(-60,345){7}
//: {8}(127,78)(127,121)(141,121){9}
input b1;    //: /sn:0 {0}(141,81)(125,81)(125,81)(114,81){1}
//: {2}(110,81)(19,81)(19,81)(-53,81){3}
//: {4}(-57,81)(-100,81)(-100,81)(-123,81){5}
//: {6}(-55,83)(-55,345){7}
//: {8}(112,83)(112,126)(141,126){9}
input a0;    //: /sn:0 {0}(141,8)(133,8)(133,8)(127,8){1}
//: {2}(123,8)(-104,8){3}
//: {4}(-108,8)(-125,8){5}
//: {6}(-106,10)(-106,344){7}
//: {8}(125,10)(125,31)(141,31){9}
input b0;    //: /sn:0 {0}(141,13)(125,13)(125,13)(112,13){1}
//: {2}(108,13)(-99,13){3}
//: {4}(-103,13)(-125,13){5}
//: {6}(-101,15)(-101,344){7}
//: {8}(110,15)(110,36)(141,36){9}
input cin;    //: /sn:0 {0}(448,69)(406,69)(406,-11){1}
//: {2}(408,-13)(444,-13)(444,6)(448,6){3}
//: {4}(404,-13)(359,-13){5}
//: {6}(355,-13)(285,-13){7}
//: {8}(281,-13)(-109,-13){9}
//: {10}(-113,-13)(-117,-13)(-117,-13)(-126,-13){11}
//: {12}(-111,-11)(-111,344){13}
//: {14}(283,-11)(283,239)(449,239){15}
//: {16}(357,-11)(357,142)(448,142){17}
output cout;    //: /sn:0 {0}(75,376)(75,360)(580,360)(580,334)(552,334){1}
wire w6;    //: /sn:0 {0}(531,34)(463,34)(463,34)(392,34){1}
//: {2}(388,34)(332,34){3}
//: {4}(328,34)(253,34){5}
//: {6}(249,34)(162,34){7}
//: {8}(251,36)(251,274)(449,274){9}
//: {10}(330,36)(330,170)(448,170){11}
//: {12}(390,36)(390,100)(447,100){13}
wire w16;    //: /sn:0 {0}(469,175)(488,175)(488,204)(533,204){1}
wire w13;    //: /sn:0 {0}(470,281)(491,281)(491,329)(531,329){1}
wire w7;    //: /sn:0 {0}(469,74)(495,74)(495,114)(531,114){1}
wire w4;    //: /sn:0 {0}(531,344)(310,344)(310,344)(160,344){1}
wire w25;    //: /sn:0 {0}(470,331)(482,331)(482,339)(531,339){1}
wire w3;    //: /sn:0 {0}(160,214)(180,214)(180,214)(201,214){1}
//: {2}(205,214)(533,214){3}
//: {4}(203,216)(203,328)(449,328){5}
wire w0;    //: /sn:0 {0}(470,249)(497,249)(497,324)(531,324){1}
wire w12;    //: /sn:0 {0}(449,313)(211,313)(211,261){1}
//: {2}(213,259)(229,259){3}
//: {4}(233,259)(449,259){5}
//: {6}(231,261)(231,289)(449,289){7}
//: {8}(209,259)(197,259){9}
//: {10}(193,259)(162,259){11}
//: {12}(195,261)(195,333)(449,333){13}
wire w18;    //: /sn:0 {0}(554,206)(564,206)(564,230)(30,230)(30,345){1}
wire w10;    //: /sn:0 {0}(-65,345)(-65,57)(575,57)(575,32)(552,32){1}
wire w24;    //: /sn:0 {0}(531,334)(485,334)(485,308)(470,308){1}
wire w1;    //: /sn:0 {0}(531,29)(504,29)(504,9)(469,9){1}
wire w8;    //: /sn:0 {0}(468,103)(487,103)(487,119)(531,119){1}
wire w17;    //: /sn:0 {0}(533,209)(485,209)(485,197)(469,197){1}
wire w14;    //: /sn:0 {0}(449,249)(268,249)(268,81){1}
//: {2}(270,79)(319,79){3}
//: {4}(323,79)(339,79){5}
//: {6}(343,79)(382,79){7}
//: {8}(386,79)(419,79)(419,79)(448,79){9}
//: {10}(384,81)(384,105)(447,105){11}
//: {12}(341,81)(341,152)(448,152){13}
//: {14}(321,81)(321,175)(448,175){15}
//: {16}(266,79)(245,79){17}
//: {18}(241,79)(199,79)(199,79)(162,79){19}
//: {20}(243,81)(243,279)(449,279){21}
wire w11;    //: /sn:0 {0}(449,284)(236,284)(236,159){1}
//: {2}(238,157)(258,157){3}
//: {4}(262,157)(289,157){5}
//: {6}(293,157)(311,157){7}
//: {8}(315,157)(382,157)(382,157)(448,157){9}
//: {10}(313,159)(313,180)(448,180){11}
//: {12}(291,159)(291,199)(448,199){13}
//: {14}(260,159)(260,254)(449,254){15}
//: {16}(234,157)(220,157){17}
//: {18}(216,157)(163,157){19}
//: {20}(218,159)(218,308)(449,308){21}
wire w2;    //: /sn:0 {0}(162,124)(191,124)(191,124)(224,124){1}
//: {2}(228,124)(297,124){3}
//: {4}(301,124)(413,124)(413,124)(531,124){5}
//: {6}(299,126)(299,194)(448,194){7}
//: {8}(226,126)(226,303)(449,303){9}
wire w15;    //: /sn:0 {0}(533,199)(496,199)(496,149)(469,149){1}
wire w5;    //: /sn:0 {0}(162,11)(217,11)(217,11)(274,11){1}
//: {2}(278,11)(347,11){3}
//: {4}(351,11)(397,11){5}
//: {6}(401,11)(427,11)(427,11)(448,11){7}
//: {8}(399,13)(399,74)(448,74){9}
//: {10}(349,13)(349,147)(448,147){11}
//: {12}(276,13)(276,244)(449,244){13}
wire w9;    //: /sn:0 {0}(552,119)(585,119)(585,134)(-21,134)(-21,346){1}
//: enddecls

  //: comment g44 @(166,144) /sn:0
  //: /line:"P2"
  //: /end
  //: IN g4 (b0) @(-127,13) /sn:0 /w:[ 5 ]
  //: comment g8 @(165,21) /sn:0
  //: /line:"G0"
  //: /end
  _GGAND3 #(8) g75 (.I0(w2), .I1(w11), .I2(w12), .Z(w24));   //: @(460,308) /sn:0 /w:[ 9 21 0 1 ]
  //: joint g47 (a3) @(123, 256) /w:[ 4 -1 3 6 ]
  //: IN g3 (cin) @(-128,-13) /sn:0 /w:[ 11 ]
  //: joint g16 (b1) @(112, 81) /w:[ 1 -1 2 8 ]
  //: joint g90 (a3) @(35, 256) /w:[ 2 -1 1 8 ]
  //: comment g17 @(167,66) /sn:0
  //: /line:"P1"
  //: /end
  _GGAND3 #(8) g26 (.I0(cin), .I1(w5), .I2(w14), .Z(w7));   //: @(459,74) /sn:0 /w:[ 0 9 9 0 ]
  //: IN g2 (a0) @(-127,8) /sn:0 /w:[ 5 ]
  //: OUT g91 (cout) @(75,373) /sn:0 /R:3 /w:[ 0 ]
  //: joint g30 (w14) @(384, 79) /w:[ 8 -1 7 10 ]
  //: joint g23 (a0) @(-106, 8) /w:[ 3 -1 4 6 ]
  //: joint g74 (w12) @(231, 259) /w:[ 4 -1 3 6 ]
  //: comment g92 @(611,202) /sn:0
  //: /line:"Count2=cin3"
  //: /end
  //: joint g86 (a2) @(-16, 154) /w:[ 2 -1 8 1 ]
  //: IN g39 (a2) @(-128,154) /sn:0 /w:[ 9 ]
  _GGOR2 #(6) g1 (.I0(a0), .I1(b0), .Z(w5));   //: @(152,11) /sn:0 /w:[ 0 0 0 ]
  //: joint g24 (b0) @(-101, 13) /w:[ 3 -1 4 6 ]
  //: joint g77 (w11) @(218, 157) /w:[ 17 -1 18 20 ]
  //: joint g29 (w6) @(390, 34) /w:[ 1 -1 2 12 ]
  //: joint g60 (w11) @(313, 157) /w:[ 8 -1 7 10 ]
  //: joint g51 (b3) @(108, 261) /w:[ 4 -1 3 6 ]
  //: joint g18 (a1) @(127, 76) /w:[ 1 -1 2 8 ]
  _GGAND4 #(10) g70 (.I0(w6), .I1(w14), .I2(w11), .I3(w12), .Z(w13));   //: @(460,281) /sn:0 /w:[ 9 21 0 7 0 ]
  _GGOR5 #(12) g82 (.I0(w0), .I1(w13), .I2(w24), .I3(w25), .I4(w4), .Z(cout));   //: @(542,334) /sn:0 /w:[ 1 1 0 1 0 1 ]
  _GGOR2 #(6) g25 (.I0(w1), .I1(w6), .Z(w10));   //: @(542,32) /sn:0 /w:[ 0 0 1 ]
  //: joint g10 (cin) @(406, -13) /w:[ 2 -1 4 1 ]
  _GGAND5 #(12) g65 (.I0(cin), .I1(w5), .I2(w14), .I3(w11), .I4(w12), .Z(w0));   //: @(460,249) /sn:0 /w:[ 15 13 0 15 5 0 ]
  _GGOR4 #(10) g64 (.I0(w15), .I1(w16), .I2(w17), .I3(w3), .Z(w18));   //: @(544,206) /sn:0 /w:[ 0 1 0 3 0 ]
  _GGAND2 #(6) g49 (.I0(a3), .I1(b3), .Z(w4));   //: @(150,344) /sn:0 /w:[ 7 7 1 ]
  //: joint g72 (w14) @(243, 79) /w:[ 17 -1 18 20 ]
  //: IN g50 (b3) @(-129,261) /sn:0 /w:[ 0 ]
  //: joint g6 (b0) @(110, 13) /w:[ 1 -1 2 8 ]
  //: joint g35 (a1) @(-60, 76) /w:[ 3 -1 4 6 ]
  //: comment g7 @(165,-2) /sn:0
  //: /line:"P0"
  //: /end
  _GGAND2 #(6) g9 (.I0(cin), .I1(w5), .Z(w1));   //: @(459,9) /sn:0 /w:[ 3 7 1 ]
  //: joint g56 (cin) @(357, -13) /w:[ 5 -1 6 16 ]
  //: joint g58 (w6) @(330, 34) /w:[ 3 -1 4 10 ]
  //: joint g68 (w14) @(268, 79) /w:[ 2 -1 16 1 ]
  //: joint g73 (w11) @(236, 157) /w:[ 2 -1 16 1 ]
  _GGOR3 #(8) g31 (.I0(w7), .I1(w8), .I2(w2), .Z(w9));   //: @(542,119) /sn:0 /w:[ 1 1 5 0 ]
  //: joint g22 (cin) @(-111, -13) /w:[ 9 -1 10 12 ]
  //: joint g59 (w14) @(321, 79) /w:[ 4 -1 3 14 ]
  //: joint g71 (w6) @(251, 34) /w:[ 5 -1 6 8 ]
  _GGXOR3 #(11) g87 (.I0(b3), .I1(a3), .I2(w18), .Z(s3));   //: @(35,356) /sn:0 /R:3 /w:[ 9 9 1 1 ]
  //: joint g85 (b2) @(-11, 159) /w:[ 2 -1 1 8 ]
  //: joint g67 (w5) @(276, 11) /w:[ 2 -1 1 12 ]
  _GGXOR3 #(11) g83 (.I0(b2), .I1(a2), .I2(w9), .Z(s2));   //: @(-16,357) /sn:0 /R:3 /w:[ 9 0 1 1 ]
  //: IN g41 (a3) @(-129,256) /sn:0 /w:[ 0 ]
  //: joint g45 (a2) @(124, 154) /w:[ 4 -1 3 6 ]
  //: joint g36 (b1) @(-55, 81) /w:[ 3 -1 4 6 ]
  _GGXOR3 #(11) g33 (.I0(b1), .I1(a1), .I2(w10), .Z(s1));   //: @(-60,356) /sn:0 /R:3 /w:[ 7 7 0 0 ]
  //: joint g54 (w14) @(341, 79) /w:[ 6 -1 5 12 ]
  //: comment g52 @(163,328) /sn:0
  //: /line:"G3"
  //: /end
  //: comment g40 @(165,244) /sn:0
  //: /line:"P3"
  //: /end
  _GGOR2 #(6) g42 (.I0(a2), .I1(b2), .Z(w11));   //: @(153,157) /sn:0 /w:[ 5 5 19 ]
  //: joint g69 (w11) @(260, 157) /w:[ 4 -1 3 14 ]
  //: joint g81 (w12) @(195, 259) /w:[ 9 -1 10 12 ]
  //: joint g66 (cin) @(283, -13) /w:[ 7 -1 8 14 ]
  //: IN g12 (b1) @(-125,81) /sn:0 /w:[ 5 ]
  _GGAND2 #(6) g46 (.I0(a2), .I1(b2), .Z(w3));   //: @(150,214) /sn:0 /w:[ 7 7 0 ]
  //: OUT g34 (s1) @(-60,373) /sn:0 /R:3 /w:[ 1 ]
  _GGAND2 #(6) g28 (.I0(w6), .I1(w14), .Z(w8));   //: @(458,103) /sn:0 /w:[ 13 11 0 ]
  _GGAND3 #(8) g57 (.I0(w6), .I1(w14), .I2(w11), .Z(w16));   //: @(459,175) /sn:0 /w:[ 11 15 11 0 ]
  //: OUT g84 (s2) @(-16,373) /sn:0 /R:3 /w:[ 0 ]
  //: joint g5 (a0) @(125, 8) /w:[ 1 -1 2 8 ]
  //: comment g11 @(608,26) /sn:0
  //: /line:"Cout0=cin1"
  //: /end
  //: IN g14 (a1) @(-125,76) /sn:0 /w:[ 5 ]
  _GGAND2 #(6) g19 (.I0(a1), .I1(b1), .Z(w2));   //: @(152,124) /sn:0 /w:[ 9 9 0 ]
  //: OUT g21 (s0) @(-106,373) /sn:0 /R:3 /w:[ 0 ]
  _GGAND2 #(6) g61 (.I0(w2), .I1(w11), .Z(w17));   //: @(459,197) /sn:0 /w:[ 7 13 1 ]
  //: comment g32 @(609,113) /sn:0
  //: /line:"Count1=cin2"
  //: /end
  _GGXOR3 #(11) g20 (.I0(b0), .I1(a0), .I2(cin), .Z(s0));   //: @(-106,355) /sn:0 /R:3 /w:[ 7 7 13 1 ]
  //: joint g78 (w12) @(211, 259) /w:[ 2 -1 8 1 ]
  _GGAND2 #(6) g79 (.I0(w3), .I1(w12), .Z(w25));   //: @(460,331) /sn:0 /w:[ 5 13 0 ]
  //: joint g63 (w11) @(291, 157) /w:[ 6 -1 5 12 ]
  //: comment g93 @(591,328) /sn:0
  //: /line:"Count3=final carry out"
  //: /end
  //: joint g89 (b3) @(40, 261) /w:[ 2 -1 1 8 ]
  //: joint g43 (b2) @(109, 159) /w:[ 4 -1 3 6 ]
  //: IN g38 (b2) @(-128,159) /sn:0 /w:[ 0 ]
  _GGAND2 #(6) g0 (.I0(a0), .I1(b0), .Z(w6));   //: @(152,34) /sn:0 /w:[ 9 9 7 ]
  _GGOR2 #(6) g15 (.I0(a1), .I1(b1), .Z(w14));   //: @(152,79) /sn:0 /w:[ 0 0 19 ]
  _GGOR2 #(6) g48 (.I0(a3), .I1(b3), .Z(w12));   //: @(152,259) /sn:0 /w:[ 5 5 11 ]
  //: joint g27 (w5) @(399, 11) /w:[ 6 -1 5 8 ]
  //: comment g37 @(165,199) /sn:0
  //: /line:"G2"
  //: /end
  //: joint g62 (w2) @(299, 124) /w:[ 4 -1 3 6 ]
  //: OUT g88 (s3) @(35,373) /sn:0 /R:3 /w:[ 0 ]
  //: joint g55 (w5) @(349, 11) /w:[ 4 -1 3 10 ]
  //: joint g80 (w3) @(203, 214) /w:[ 2 -1 1 4 ]
  //: comment g13 @(167,111) /sn:0
  //: /line:"G1"
  //: /end
  _GGAND4 #(10) g53 (.I0(cin), .I1(w5), .I2(w14), .I3(w11), .Z(w15));   //: @(459,149) /sn:0 /w:[ 17 11 13 9 1 ]
  //: joint g76 (w2) @(226, 124) /w:[ 2 -1 1 8 ]

endmodule
//: /netlistEnd

