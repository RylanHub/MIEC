//: version "2.1"
//: property encoding = "utf-8"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "Lab5_A.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
supply1 w6;    //: /sn:0 {0}(267,173)(174,173){1}
//: {2}(172,171)(172,105){3}
//: {4}(172,175)(172,239)(267,239){5}
reg w1;    //: /sn:0 {0}(267,205)(236,205)(236,315){1}
//: {2}(238,317)(474,317)(474,215)(574,215){3}
//: {4}(234,317)(201,317){5}
reg w2;    //: /sn:0 {0}(641,283)(641,337)(336,337){1}
//: {2}(334,335)(334,273){3}
//: {4}(334,339)(334,354){5}
wire w4;    //: /sn:0 {0}(404,224)(419,224){1}
wire [1:0] w3;    //: /sn:0 {0}(#:466,132)(466,113){1}
wire w10;    //: /sn:0 {0}(711,234)(726,234){1}
wire w5;    //: /sn:0 {0}(574,183)(510,183){1}
//: {2}(506,183)(473,183){3}
//: {4}(471,181)(471,138){5}
//: {6}(469,183)(404,183){7}
//: {8}(508,185)(508,249)(574,249){9}
wire w9;    //: /sn:0 {0}(461,138)(461,153)(737,153)(737,193)(711,193){1}
//: enddecls

  //: LED g8 (w3) @(466,106) /sn:0 /w:[ 1 ] /type:3
  //: joint g4 (w5) @(508, 183) /w:[ 1 -1 2 8 ]
  //: SWITCH g3 (w1) @(184,317) /sn:0 /w:[ 5 ] /st:0 /dn:0
  //: joint g2 (w6) @(172, 173) /w:[ 1 2 -1 4 ]
  //: VDD g1 (w6) @(183,105) /sn:0 /w:[ 3 ]
  //: joint g10 (w5) @(471, 183) /w:[ 3 4 6 -1 ]
  //: SWITCH g6 (w2) @(334,368) /sn:0 /R:1 /w:[ 5 ] /st:0 /dn:0
  assign w3 = {w9, w5}; //: CONCAT g9  @(466,133) /sn:0 /R:1 /w:[ 0 0 5 ] /dr:0 /tp:0 /drp:1
  //: joint g7 (w2) @(334, 337) /w:[ 1 2 -1 4 ]
  //: joint g11 (w1) @(236, 317) /w:[ 2 1 4 -1 ]
  JKFlipFlop g5 (.J(w5), .K(w5), .CLOCK(w1), .RESET(w2), .Q(w9), .Qinv(w10));   //: @(575, 164) /sz:(135, 118) /sn:0 /p:[ Li0>0 Li1>9 Li2>3 Bi0>0 Ro0<1 Ro1<0 ]
  JKFlipFlop g0 (.J(w6), .K(w6), .CLOCK(w1), .RESET(w2), .Q(w5), .Qinv(w4));   //: @(268, 154) /sz:(135, 118) /sn:0 /p:[ Li0>0 Li1>5 Li2>0 Bi0>3 Ro0<7 Ro1<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin JKFlipFlop
module JKFlipFlop(CLOCK, RESET, Q, K, Qinv, J);
//: interface  /sz:(135, 118) /bd:[ Li0>CLOCK(51/118) Li1>K(85/118) Li2>J(19/118) Bi0>RESET(66/135) Ro0<Qinv(70/118) Ro1<Q(29/118) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input CLOCK;    //: /sn:0 {0}(256,222)(240,222)(240,253){1}
//: {2}(238,255)(227,255)(227,348){3}
//: {4}(229,350)(242,350){5}
//: {6}(246,350)(256,350){7}
//: {8}(244,352)(244,355)(256,355){9}
//: {10}(225,350)(205,350){11}
//: {12}(240,257)(240,288)(255,288){13}
output Q;    //: /sn:0 {0}(642,226)(578,226)(578,226)(602,226){1}
//: {2}(598,226)(542,226){3}
//: {4}(538,226)(524,226){5}
//: {6}(540,228)(540,258)(486,258)(486,286)(506,286){7}
//: {8}(600,228)(600,330)(242,330)(242,298)(255,298){9}
input K;    //: /sn:0 {0}(255,293)(239,293)(239,293)(204,293){1}
input RESET;    //: /sn:0 {0}(382,380)(382,321){1}
//: {2}(384,319)(491,319)(491,296)(506,296){3}
//: {4}(380,319)(331,319)(331,298)(346,298){5}
input J;    //: /sn:0 {0}(256,217)(241,217)(241,217)(208,217){1}
output Qinv;    //: /sn:0 {0}(640,291)(609,291)(609,291)(588,291){1}
//: {2}(586,289)(586,177)(230,177)(230,212)(256,212){3}
//: {4}(584,291)(571,291){5}
//: {6}(569,289)(569,251)(494,251)(494,228)(503,228){7}
//: {8}(567,291)(564,291)(564,291)(527,291){9}
wire w6;    //: /sn:0 {0}(346,293)(330,293)(330,293)(276,293){1}
wire w7;    //: /sn:0 {0}(458,293)(443,293)(443,293)(393,293){1}
//: {2}(391,291)(391,255)(328,255)(328,222)(352,222){3}
//: {4}(389,293)(367,293){5}
wire w4;    //: /sn:0 {0}(451,220)(430,220)(430,220)(387,220){1}
//: {2}(383,220)(373,220){3}
//: {4}(385,222)(385,262)(319,262)(319,288)(346,288){5}
wire w14;    //: /sn:0 {0}(479,291)(494,291)(494,291)(506,291){1}
wire w2;    //: /sn:0 {0}(352,217)(303,217)(303,217)(277,217){1}
wire w5;    //: /sn:0 {0}(503,223)(488,223)(488,223)(472,223){1}
wire w9;    //: /sn:0 {0}(458,288)(438,288)(438,257){1}
//: {2}(438,253)(438,225)(451,225){3}
//: {4}(436,255)(420,255)(420,353)(277,353){5}
//: enddecls

  //: joint g8 (CLOCK) @(244, 350) /w:[ 6 -1 5 8 ]
  _GGNAND3 #(6) g4 (.I0(CLOCK), .I1(K), .I2(Q), .Z(w6));   //: @(266,293) /sn:0 /w:[ 13 0 9 1 ]
  _GGNAND3 #(6) g16 (.I0(Q), .I1(w14), .I2(RESET), .Z(Qinv));   //: @(517,291) /sn:0 /w:[ 7 1 3 9 ]
  _GGNAND3 #(6) g3 (.I0(Qinv), .I1(J), .I2(CLOCK), .Z(w2));   //: @(267,217) /sn:0 /w:[ 3 0 0 1 ]
  //: joint g17 (Q) @(540, 226) /w:[ 3 -1 4 6 ]
  //: IN g2 (CLOCK) @(203,350) /sn:0 /w:[ 11 ]
  //: IN g23 (RESET) @(382,382) /sn:0 /R:1 /w:[ 0 ]
  //: OUT g24 (Q) @(639,226) /sn:0 /w:[ 0 ]
  //: IN g1 (K) @(202,293) /sn:0 /w:[ 1 ]
  //: joint g18 (Qinv) @(569, 291) /w:[ 5 6 8 -1 ]
  //: OUT g25 (Qinv) @(637,291) /sn:0 /w:[ 0 ]
  //: joint g10 (CLOCK) @(227, 350) /w:[ 4 3 10 -1 ]
  _GGNAND2 #(4) g6 (.I0(w2), .I1(w7), .Z(w4));   //: @(363,220) /sn:0 /w:[ 0 3 3 ]
  //: joint g9 (CLOCK) @(240, 255) /w:[ -1 1 2 12 ]
  _GGNAND3 #(6) g7 (.I0(w4), .I1(w6), .I2(RESET), .Z(w7));   //: @(357,293) /sn:0 /w:[ 5 0 5 5 ]
  //: joint g22 (Q) @(600, 226) /w:[ 1 -1 2 8 ]
  //: joint g12 (w4) @(385, 220) /w:[ 1 -1 2 4 ]
  _GGNAND2 #(4) g14 (.I0(w5), .I1(Qinv), .Z(Q));   //: @(514,226) /sn:0 /w:[ 0 7 5 ]
  //: joint g11 (w7) @(391, 293) /w:[ 1 2 4 -1 ]
  _GGNAND2 #(4) g5 (.I0(CLOCK), .I1(CLOCK), .Z(w9));   //: @(267,353) /sn:0 /w:[ 7 9 5 ]
  //: joint g19 (RESET) @(382, 319) /w:[ 2 -1 4 1 ]
  //: joint g21 (Qinv) @(586, 291) /w:[ 1 2 4 -1 ]
  //: joint g20 (w9) @(438, 255) /w:[ -1 2 4 1 ]
  _GGNAND2 #(4) g15 (.I0(w9), .I1(w7), .Z(w14));   //: @(469,291) /sn:0 /w:[ 0 0 0 ]
  //: IN g0 (J) @(206,217) /sn:0 /w:[ 1 ]
  _GGNAND2 #(4) g13 (.I0(w4), .I1(w9), .Z(w5));   //: @(462,223) /sn:0 /w:[ 0 3 1 ]

endmodule
//: /netlistEnd

