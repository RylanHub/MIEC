//: version "2.1"
//: property encoding = "utf-8"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "Lab3.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg A0;    //: /sn:0 {0}(172,113)(311,113){1}
//: {2}(315,113)(357,113)(357,140)(368,140){3}
//: {4}(313,115)(313,233)(371,233){5}
reg B1;    //: /sn:0 {0}(271,465)(183,465){1}
reg A1;    //: /sn:0 {0}(181,420)(320,420){1}
//: {2}(324,420)(366,420)(366,447)(377,447){3}
//: {4}(322,422)(322,540)(380,540){5}
reg S;    //: /sn:0 {0}(99,303)(139,303){1}
//: {2}(143,303)(481,303)(481,221){3}
//: {4}(483,219)(610,219){5}
//: {6}(481,217)(481,177)(612,177){7}
//: {8}(141,301)(141,258)(228,258){9}
//: {10}(230,256)(230,163)(248,163){11}
//: {12}(230,260)(230,470)(271,470){13}
reg B0;    //: /sn:0 {0}(248,158)(174,158){1}
wire w6;    //: /sn:0 {0}(392,236)(673,236){1}
wire w7;    //: /sn:0 {0}(647,159)(647,175)(633,175){1}
wire w4;    //: /sn:0 {0}(612,172)(581,172)(581,143)(548,143){1}
//: {2}(544,143)(389,143){3}
//: {4}(546,145)(546,214)(610,214){5}
wire w10;    //: /sn:0 {0}(673,231)(659,231)(659,217)(631,217){1}
wire w8;    //: /sn:0 {0}(656,466)(656,483)(650,483){1}
wire w14;    //: /sn:0 {0}(704,511)(704,541)(703,541){1}
wire Z1;    //: /sn:0 {0}(694,234)(749,234)(749,387)(476,387)(476,507)(492,507){1}
//: {2}(494,505)(494,485)(629,485){3}
//: {4}(494,509)(494,526)(619,526){5}
wire w11;    //: /sn:0 {0}(682,538)(668,538)(668,524)(640,524){1}
wire w5;    //: /sn:0 {0}(629,480)(598,480)(598,450)(557,450){1}
//: {2}(553,450)(398,450){3}
//: {4}(555,452)(555,521)(619,521){5}
wire Y0;    //: /sn:0 {0}(269,161)(297,161){1}
//: {2}(301,161)(355,161)(355,145)(368,145){3}
//: {4}(299,163)(299,238)(371,238){5}
wire w9;    //: /sn:0 {0}(401,543)(682,543){1}
wire Y1;    //: /sn:0 {0}(292,468)(306,468){1}
//: {2}(310,468)(364,468)(364,452)(377,452){3}
//: {4}(308,470)(308,545)(380,545){5}
//: enddecls

  _GGXOR2 #(8) g8 (.I0(w5), .I1(Z1), .Z(w8));   //: @(640,483) /sn:0 /w:[ 0 3 1 ]
  //: SWITCH g4 (A1) @(164,420) /sn:0 /w:[ 0 ] /st:1 /dn:1
  //: SWITCH A0 (A0) @(155,113) /sn:0 /w:[ 0 ] /st:1 /dn:1
  //: LED S1 (w8) @(656,459) /w:[ 0 ] /type:0
  //: joint g3 (A0) @(313, 113) /w:[ 2 -1 1 4 ]
  //: joint g16 (w4) @(546, 143) /w:[ 1 -1 2 4 ]
  _GGXOR2 #(8) g17 (.I0(w4), .I1(S), .Z(w7));   //: @(623,175) /sn:0 /w:[ 0 7 1 ]
  //: joint g2 (Y0) @(299, 161) /w:[ 2 -1 1 4 ]
  _GGAND2 #(6) g23 (.I0(A1), .I1(Y1), .Z(w9));   //: @(391,543) /sn:0 /w:[ 5 5 0 ]
  _GGOR2 #(6) g24 (.I0(w11), .I1(w9), .Z(w14));   //: @(693,541) /sn:0 /w:[ 0 1 1 ]
  _GGXOR2 #(8) g1 (.I0(B0), .I1(S), .Z(Y0));   //: @(259,161) /sn:0 /w:[ 0 11 0 ]
  //: SWITCH g18 (S) @(82,303) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: joint g25 (S) @(230, 258) /w:[ -1 10 9 12 ]
  _GGXOR2 #(8) g10 (.I0(B1), .I1(S), .Z(Y1));   //: @(282,468) /sn:0 /w:[ 0 13 0 ]
  //: joint g6 (w5) @(555, 450) /w:[ 1 -1 2 4 ]
  //: joint g9 (Y1) @(308, 468) /w:[ 2 -1 1 4 ]
  //: joint g7 (A1) @(322, 420) /w:[ 2 -1 1 4 ]
  _GGXOR2 #(8) g22 (.I0(A0), .I1(Y0), .Z(w4));   //: @(379,143) /sn:0 /w:[ 3 3 3 ]
  //: LED C2 (w14) @(704,504) /w:[ 0 ] /type:0
  //: LED S0 (w7) @(647,152) /w:[ 0 ] /type:0
  _GGXOR2 #(8) g12 (.I0(A1), .I1(Y1), .Z(w5));   //: @(388,450) /sn:0 /w:[ 3 3 3 ]
  //: SWITCH g28 (B1) @(166,465) /sn:0 /w:[ 1 ] /st:0 /dn:1
  _GGAND2 #(6) g14 (.I0(A0), .I1(Y0), .Z(w6));   //: @(382,236) /sn:0 /w:[ 5 5 0 ]
  _GGAND2 #(6) g5 (.I0(w4), .I1(S), .Z(w10));   //: @(621,217) /sn:0 /w:[ 5 5 1 ]
  //: joint g21 (S) @(141, 303) /w:[ 2 8 1 -1 ]
  _GGOR2 #(6) g19 (.I0(w10), .I1(w6), .Z(Z1));   //: @(684,234) /sn:0 /w:[ 0 1 0 ]
  //: joint g20 (S) @(481, 219) /w:[ 4 6 -1 3 ]
  //: joint g15 (Z1) @(494, 507) /w:[ -1 2 1 4 ]
  //: SWITCH g0 (B0) @(157,158) /sn:0 /w:[ 1 ] /st:1 /dn:1
  _GGAND2 #(6) g13 (.I0(w5), .I1(Z1), .Z(w11));   //: @(630,524) /sn:0 /w:[ 5 5 1 ]

endmodule
//: /netlistEnd

